** Profile: "SCHEMATIC1-Circuit"  [ C:\Users\zobay\OneDrive\Desktop\Thesis defense\TCAM circuit\tcam -pspicefiles\schematic1\circuit.sim ] 

** Creating circuit file "Circuit.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Cadence/SPB_16.6/tools/capture/library/pspice/memristor.lib" 
* From [PSPICE NETLIST] section of C:\Users\zobay\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 200ms 0 
.OPTIONS ADVCONV
.OPTIONS DIGINITSTATE= 0
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
